module random(
    input CLK // Clock
    , output[7:0] DAT_OUT // Output random number
    , input ASYNC_RST_L // Async reset (low-level)
);
endmodule
